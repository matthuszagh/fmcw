`define FMCW_PARAMS parameter \
GPIO_WIDTH = 6, \
USB_DATA_WIDTH = 8, \
ADC_DATA_WIDTH = 12, \
SD_DATA_WIDTH = 4, \
FIR_M = 20, \
FIR_M_WIDTH = 5, \
FIR_INPUT_WIDTH = 12, \
FIR_INTERNAL_WIDTH = 39, \
FIR_NORM_SHIFT = 4, \
FIR_OUTPUT_WIDTH = 14, \
FIR_TAP_WIDTH = 16, \
FIR_POLY_BANK_LEN = 60, \
FIR_POLY_BANK_LEN_LOG2 = 6, \
FIR_ROM_SIZE = 128, \
FFT_TWIDDLE_WIDTH = 10, \
FFT_DIST_N = 1024, \
FFT_DIST_N_LOG2 = 10, \
FFT_DIST_N_STAGES = 5, \
FFT_DIST_INPUT_WIDTH = 14, \
FFT_DIST_INTERNAL_WIDTH = 25, \
FFT_DIST_OUTPUT_WIDTH = 25, \
FFT_ANGLE_N = 256, \
FFT_ANGLE_N_LOG2 = 8, \
FFT_ANGLE_N_STAGES = 4, \
FFT_ANGLE_INPUT_WIDTH = 14, \
FFT_ANGLE_INTERNAL_WIDTH = 23, \
FFT_ANGLE_OUTPUT_WIDTH = 23