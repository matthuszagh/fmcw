`define FMCW_DEFAULT_PARAMS parameter \
NTAPS = 120, \
CntW = 7, \
TW = 16, \
IW = 12, \
OW = 16, \
IntW = 29, \
M = 20, \
MW = 5
