`define FMCW_DEFAULT_PARAMS parameter \
NTAPS = 120, \
CntW = 7, \
TW = 16, \
IW = 12, \
OW = 24, \
IntW = 29, \
USBDW = 8, \
SDDW = 4, \
GPIOW = 6, \
FFT_N = 1024, \
FFT_STAGES = 5, \
FFT_NLOG2 = 10, \
FFTDW = 32, \
TWIDDLE_WIDTH = 10, \
Cnt_STAGE = 3, \
M = 20, \
MW = 5
