`ifndef _FT245_V_
`define _FT245_V_

`default_nettype none
`timescale 1ns/1ps

/** ft245.v
 *
 * An interface for using the FT2232H chip in FT245 synchronous FIFO
 * mode.
 */

`include "async_fifo.v"
`include "pll_sync_ctr.v"

`define FT_DATA_WIDTH 8
`define CLK_FREQ 40000000
`define FLUSH_PERIOD 10  // 10 periods of 40MHz in 250ns
`define READ_SUCCESS 8'b1000_1110
`define READ_FAILURE 8'b1000_0000

module ft245 #(
   // The FIFO is used to buffer write data when the FT2232H's
   // internal buffer is full. It also prevents CDC issues since `clk'
   // and `ft_clk' are asynchronous.
   parameter WRITE_DEPTH    = 1024,
   // A FIFO used to buffer read data from FT2232H to FPGA.
   parameter READ_DEPTH     = 512,
   // The number of bits in a payload (does not include header/tail
   // and other bits). This must be less than or equal to 52. For any
   // number less than 52, the remaining bits will be set to 0. The
   // zero bits will appear as the most significant bits in the 52 bit
   // range.
   parameter DATA_WIDTH     = 39,
   // Duplicate all transmission bytes as a form of error
   // detection. Although inefficient, this is effective at avoiding
   // data errors caused by the host PC missing bytes while reading.
   parameter DUPLICATE_TX   = 1
) (
   // ======================== FPGA interface ========================

   // A reset signal is required to start the FIFO in a known state.
   input wire                      rst_n,
   // Synchronizes reads and writes between the FT245 and FPGA. This
   // clock does not require any known phase relation to `ft_clk'.
   input wire                      clk,
   // Pull high to write data from FPGA to FT2232H for transmission to
   // host PC.
   input wire                      wren,
   // Write data.
   input wire [DATA_WIDTH-1:0]     wrdata,
   output wire                     wrfifo_full,
   output wire                     wrfifo_empty,
   // Pull high to read data from internal read FIFO. It only makes
   // sense to read data when !rdfifo_empty.
   input wire                      rden,
   output reg [DATA_WIDTH-1:0]     rddata,
   output wire                     rdfifo_full,
   output wire                     rdfifo_empty,

   // ========================= PC interface =========================

   // Most of these ports should be connected directly to the
   // corresponding IO ports on the FPGA.

   // Clock generated by the FT2232H and used to synchronize data
   // transfers.
   input wire                      ft_clk,
   // Synchronizes write word changes. `slow_ft_clk' * `DATA_WIDTH' /
   // 8 = `ft_clk'.
   input wire                      slow_ft_clk,
   // Low indicates there is data available to be read from the FIFO.
   input wire                      rxf_n,
   // Low indicates data can be written to the FIFO.
   input wire                      txe_n,
   // 0 makes read data from the FIFO available at the data pins.
   output reg                      rd_n,
   // Pull low to register write data from the data pins into the
   // FIFO.
   output reg                      wr_n,
   // Drive low to read data from FIFO. Must be deasserted at least 1
   // clock period (`ft_clk') before driving `rd_n' low.
   output reg                      oe_n,
   // Low when USB in suspend mode.
   /* verilator lint_off UNUSED */
   input wire                      suspend_n,
   /* verilator lint_on UNUSED */
   // Strobing low (min 250ns) sends FIFO data immediately to the host
   // PC.
   output reg                      ft_siwua_n,
   inout wire [`FT_DATA_WIDTH-1:0] ft_data
);

   // TODO should be present but not supported by vivado.
   // assert (DATA_WIDTH <= 52)
   //   else $error("FT245 DATA_WIDTH must be no greater than 52 bits.");

   // number of bits in full transmission, including header/tail/meta
   // data.
   localparam FULL_WIDTH     = 64;
   localparam NBYTES         = FULL_WIDTH/8;
   localparam LEADING_BLANKS = 52 - DATA_WIDTH;
   localparam CTR_WIDTH = $clog2(NBYTES);

   // TODO this should be parameterized to work with different word
   // sizes.
`ifndef __ICARUS__
   if (NBYTES != 8) $error();
`endif

   wire [`FT_DATA_WIDTH-1:0]       rdfifo_rddata;
   wire                            rdfifo_rden;

   // Read FIFO
   async_fifo #(
     .WIDTH (`FT_DATA_WIDTH ),
     .SIZE  (READ_DEPTH     )
   ) fifo_read (
      .rst_n  (rst_n         ),
      .full   (rdfifo_full   ),
      .empty  (rdfifo_empty  ),
      .rdclk  (clk           ),
      .rden   (rdfifo_rden   ),
      .rddata (rdfifo_rddata ),
      .wrclk  (ft_clk        ),
      .wren   (!rd_n         ),
      .wrdata (ft_data       )
   );

   assign ft_data = oe_n ? ft_data_reg : 8'bzzzz_zzzz;

   wire [DATA_WIDTH-1:0]        wrfifo_rddata;
   reg [DATA_WIDTH-1:0]         wrfifo_wrdata;
   wire                         wrfifo_rden;
   // Write FIFO
   /* verilator lint_off PINMISSING */
   async_fifo #(
      .WIDTH (DATA_WIDTH  ),
      .SIZE  (WRITE_DEPTH )
   ) fifo_write (
      .rst_n  (rst_n                         ),
      .full   (wrfifo_full                   ),
      .empty  (wrfifo_empty                  ),
      .rdclk  (slow_ft_clk                   ),
      // txe_n is a guard against writes to a full buffer, since
      // FT2232H can take up to 7.15ns to report a full buffer.
      .rden   (oe_n && wrfifo_rden && !txe_n ),
      .rddata (wrfifo_rddata                 ),
      .wrclk  (clk                           ),
      .wren   (wren && !wrfifo_full          ),
      .wrdata (wrfifo_wrdata                 )
   );
   /* verilator lint_on PINMISSING */

   wire [CTR_WIDTH-1:0]         ctr;
   pll_sync_ctr #(
      .RATIO (NBYTES)
   ) pll_sync_ctr (
      .fst_clk (ft_clk      ),
      .slw_clk (slow_ft_clk ),
      .rst_n   (rst_n       ),
      .ctr     (ctr         )
   );

   reg [7:0]                    ft_data_reg;
   wire [FULL_WIDTH-1:0]        wrfifo_rddata_full;

   assign wrfifo_rddata_full = {8'h80, {LEADING_BLANKS{1'b0}}, wrfifo_rddata, 4'h0};

   always @(*) begin
      case (ctr)
      3'b000 : ft_data_reg = wrfifo_rddata_full[63:56];
      3'b001 : ft_data_reg = wrfifo_rddata_full[55:48];
      3'b010 : ft_data_reg = wrfifo_rddata_full[47:40];
      3'b011 : ft_data_reg = wrfifo_rddata_full[39:32];
      3'b100 : ft_data_reg = wrfifo_rddata_full[31:24];
      3'b101 : ft_data_reg = wrfifo_rddata_full[23:16];
      3'b110 : ft_data_reg = wrfifo_rddata_full[15:8];
      3'b111 : ft_data_reg = wrfifo_rddata_full[7:0];
      endcase
   end

   // Wait for an indication to read data from or send data to the
   // host.
   localparam [2:0] IDLE_STATE         = 3'd0;
   // Attempt to read 8 bytes from the host. If a timeout occurs
   // before 8 bytes are read, indicate a failure and request that the
   // host repeat the transmission (see ``READ_FAILURE_STATE``). If
   // the 8 bytes are read before a timeout, indicate a success (see
   // ``READ_SUCCESS_STATE``).
   localparam [2:0] READ_STATE         = 3'd1;
   // Read from host was successful. Communicate this to the host and
   // then return to idle.
   localparam [2:0] READ_SUCCESS_STATE = 3'd2;
   // Read from host failed. Communicate this to the host, requesting
   // data be repeated and then return to idle. If the host misses the
   // success or failure indication, it will assume a failure and
   // resend the transmission after a timeout.
   localparam [2:0] READ_FAILURE_STATE = 3'd3;
   // Ensure all transmission data has been received by the host
   // before proceeding.
   localparam [2:0] FLUSH_OUTPUT_STATE = 3'd4;
   // Stream data from the FPGA to the host. Stop streaming if we
   // receive data from the host.
   localparam [2:0] STREAM_STATE       = 3'd5;

   reg [2:0]                   state;
   reg [CTR_WIDTH-1:0]         rd_ctr;
   localparam [CTR_WIDTH-1:0]  RD_CTR_MAX = `FT_DATA_WIDTH - 1;
   /** Allow reads 1s before timing out. This is probably excessive,
   /* but since Linux provides no realtime guarantee, this should
   /* avoid unnecessary timeouts. */
   reg [$clog2(`CLK_FREQ)-1:0] read_timeout;
   localparam [$clog2(`CLK_FREQ)-1:0] READ_TIMEOUT_MAX = `CLK_FREQ - 1;
   reg [$clog2(`FLUSH_PERIOD)-1:0] flush_ctr;
   localparam [$clog2(`FLUSH_PERIOD)-1:0] FLUSH_CTR_MAX = `FLUSH_PERIOD - 1;
   reg                             read_status_toggle;

   always @(posedge clk) begin
      if (!rst_n) begin
         state              <= IDLE_STATE;
         rd_ctr             <= {CTR_WIDTH{1'b0}};
         read_timeout       <= {$clog2(`CLK_FREQ){1'b0}};
         flush_ctr          <= {$clog2(`FLUSH_PERIOD){1'b0}};
         read_status_toggle <= 1'b0;
      end else begin
         case (state)
         IDLE_STATE:
           begin
              if (!rdfifo_empty) begin
                 state <= READ_STATE;
              end else if (!wrfifo_empty) begin
                 state <= STREAM_STATE;
              end
              rd_ctr             <= {CTR_WIDTH{1'b0}};
              read_timeout       <= {$clog2(`CLK_FREQ){1'b0}};
              flush_ctr          <= {$clog2(`FLUSH_PERIOD){1'b0}};
              read_status_toggle <= 1'b0;
           end

         READ_STATE:
           begin
              if (!rdfifo_empty) begin
                 rddata[rd_ctr] <= rdfifo_rddata;
                 if (rd_ctr == RD_CTR_MAX) begin
                    rd_ctr       <= {CTR_WIDTH{1'b0}};
                    read_timeout <= {$clog2(`CLK_FREQ){1'b0}};
                    state        <= READ_SUCCESS_STATE;
                 end else begin
                    rd_ctr       <= rd_ctr + 1'b1;
                    read_timeout <= read_timeout + 1'b1;
                 end
              end else begin
                 if (read_timeout == READ_TIMEOUT_MAX) begin
                    rd_ctr       <= {CTR_WIDTH{1'b0}};
                    read_timeout <= {$clog2(`CLK_FREQ){1'b0}};
                    state        <= READ_FAILURE_STATE;
                 end else begin
                    read_timeout <= read_timeout + 1'b1;
                 end
              end
              flush_ctr          <= {$clog2(`FLUSH_PERIOD){1'b0}};
              read_status_toggle <= 1'b0;
           end

         READ_SUCCESS_STATE:
           begin
              if (read_status_toggle) begin
                 state <= FLUSH_OUTPUT_STATE;
              end else begin
                 wrfifo_wrdata <= `READ_SUCCESS;
              end
              rd_ctr       <= {CTR_WIDTH{1'b0}};
              read_timeout <= {$clog2(`CLK_FREQ){1'b0}};
              flush_ctr    <= {$clog2(`FLUSH_PERIOD){1'b0}};
           end

         READ_FAILURE_STATE:
           begin
              rd_ctr       <= {CTR_WIDTH{1'b0}};
              read_timeout <= {$clog2(`CLK_FREQ){1'b0}};
              flush_ctr    <= {$clog2(`FLUSH_PERIOD){1'b0}};
           end

         FLUSH_OUTPUT_STATE:
           begin
              if (flush_ctr == FLUSH_CTR_MAX) begin
                 flush_ctr <= {$clog2(`FLUSH_PERIOD){1'b0}};
                 state     <= IDLE_STATE;
              end else begin
                 flush_ctr <= flush_ctr + 1'b1;
              end
              rd_ctr       <= {CTR_WIDTH{1'b0}};
              read_timeout <= {$clog2(`CLK_FREQ){1'b0}};
           end

         STREAM_STATE:
           begin
              if (!rdfifo_empty) begin
                 state <= READ_STATE;
              end else begin
              end
              rd_ctr       <= {CTR_WIDTH{1'b0}};
              read_timeout <= {$clog2(`CLK_FREQ){1'b0}};
              flush_ctr    <= {$clog2(`FLUSH_PERIOD){1'b0}};
           end

         endcase
      end
   end

   always @(*) begin
      case (state)
      IDLE_STATE:
        begin
           rdfifo_rden = 1'b0;
           ft_siwua_n  = 1'b1;
        end

      READ_STATE:
        begin
           rdfifo_rden = 1'b1;
           ft_siwua_n  = 1'b1;
        end

      READ_SUCCESS_STATE:
        begin
           rdfifo_rden = 1'b0;
           ft_siwua_n  = 1'b1;
        end

      READ_FAILURE_STATE:
        begin
           rdfifo_rden = 1'b0;
           ft_siwua_n  = 1'b1;
        end

      FLUSH_OUTPUT_STATE:
        begin
           rdfifo_rden = 1'b0;
           ft_siwua_n  = 1'b0;
        end

      STREAM_STATE:
        begin
           rdfifo_rden = 1'b0;
           ft_siwua_n  = 1'b1;
        end

      endcase
   end


   // ================================================================




   generate
      if (DUPLICATE_TX == 1) begin
         reg duplicate;
         always @(posedge slow_ft_clk) begin
            if (!rst_n) begin
               duplicate <= 1'b0;
            end else begin
               duplicate <= ~duplicate;
            end
         end

         assign wrfifo_rden = ~duplicate;
         always @(posedge ft_clk) begin
            if (!rst_n) begin
               rd_n <= 1'b1;
               wr_n <= 1'b1;
               oe_n <= 1'b1;
               ft_siwua_n <= 1'b1;
            // favor reads
            end else if (!rxf_n) begin
               oe_n <= 1'b0;
               wr_n <= 1'b1;
               if (!oe_n) begin
                  rd_n <= 1'b0;
               end
            end else if (!txe_n) begin
               oe_n <= 1'b1;
               rd_n <= 1'b1;
               if (oe_n)
                 wr_n <= 1'b0;
            end else begin
               oe_n <= 1'b1;
               rd_n <= 1'b1;
               wr_n <= 1'b1;
            end
         end
      end else begin
         assign wrfifo_rden = 1'b1;
         always @(posedge ft_clk) begin
            if (!rst_n) begin
               rd_n <= 1'b1;
               wr_n <= 1'b1;
               oe_n <= 1'b1;
               ft_siwua_n <= 1'b1;
            end else if (!rxf_n) begin
               oe_n <= 1'b0;
               wr_n <= 1'b1;
               if (!oe_n) begin
                  rd_n <= 1'b0;
               end
            end else if (!txe_n) begin
               oe_n <= 1'b1;
               rd_n <= 1'b1;
               if (oe_n)
                 wr_n <= 1'b0;
            end else begin
               oe_n <= 1'b1;
               rd_n <= 1'b1;
               wr_n <= 1'b1;
            end
         end
      end
   endgenerate

`ifdef COCOTB_SIM
   `ifdef FT245
   initial begin
      $dumpfile ("cocotb/build/ft245.vcd");
      $dumpvars (0, ft245);
      #1;
   end
   `endif
`endif

endmodule

`undef FT_DATA_WIDTH
`undef CLK_FREQ
`undef FLUSH_PERIOD
`undef READ_SUCCESS
`undef READ_FAILURE

`endif
