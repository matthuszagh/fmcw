`default_nettype none

`include "fmcw_defines.vh"

module fft_r22sdf_rom_s0 #( `FMCW_DEFAULT_PARAMS )
   (
    input wire clk
    input wire [FFT_NLOG2-1:0] addr,
    input
    );

   initial begin

   end

endmodule // fft_r22sdf_rom_s0
